module control_unit_tb;

endmodule