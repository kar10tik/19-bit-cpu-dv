module logical_unit_tb;

endmodule