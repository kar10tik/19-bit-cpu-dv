module arithmetic_unit_tb;

endmodule