//TODO Constraints on addresses, data