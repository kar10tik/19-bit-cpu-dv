`ifndef constants_h
`define constants_h

localparam WORD_SIZE = 19;
localparam ADDR_SIZE = 20;
localparam OPCODE_SIZE = 5;

`endif