module data_memory(control_bus_if ctrl_bus_if);
    
endmodule