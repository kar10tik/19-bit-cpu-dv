module arith_logic_unit_tb;

endmodule