module data_memory_tb;

endmodule