//LUT for control signals for various opcodes
import opcodes::*;
package control_signals;

endpackage