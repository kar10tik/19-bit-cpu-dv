module register_tb;

endmodule