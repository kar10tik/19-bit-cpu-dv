module instruction_memory_tb;

endmodule